//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:   
// Design Name: 
// Module Name:    spart 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module spart(
    input clk, //Runs at 50MHz
    input rst,
    input iocs,
    input iorw,
    output rda,
    output tbr,
    input [1:0] ioaddr,
    inout [7:0] databus,
    output txd,
    input rxd
    );


    ////////////////Declared Variables//////////////////








    ////////////////Instantated Modules/////////////////







    ///////////////////////Logic///////////////////////






    //IO addressing

    //00 -> Transmit Buffer (IOR/W = 0) : Receive Buffer (IOR/W)

endmodule
